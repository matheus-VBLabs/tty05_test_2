

//IMPORTED BLOCK:bus_to_wires
// Bloco separador de barramento de 8 bits para uso na ferramenta 
module bus_to_wires (in,out_0,out_1,out_2,out_3,out_4,out_5,out_6,out_7);

// Inputs e Outputs
input wire [7:0] in;
output wire out_0,out_1,out_2,out_3,out_4,out_5,out_6,out_7;

// Comportamento do circuito
assign out_0 = in[0];
assign out_1 = in[1];
assign out_2 = in[2];
assign out_3 = in[3];
assign out_4 = in[4];
assign out_5 = in[5];
assign out_6 = in[6];
assign out_7 = in[7];

endmodule




//IMPORTED BLOCK:pulse_count_8_bits
module pulse_count_8_bits(pulse, counter);
input wire pulse;
output reg [7:0] counter;

initial counter = 0;

always @(posedge pulse) begin
counter <= counter + 1;
end

endmodule


// Automatically generated by ChipInventor Cloud EDA Tool - 2.0
// Careful: this file (hdl.v) will be automatically replaced when you ask
// to generate code from BLOCKS buttons.
module tt_um_counter_8bits (
    input  wire [7:0] ui_in,    // Dedicated inputs - connected to the input switches
    output wire [7:0] uo_out,   // Dedicated outputs - connected to the 7 segment display
    input  wire [7:0] uio_in,   // IOs: Bidirectional Input path
    output wire [7:0] uio_out,  // IOs: Bidirectional Output path
    output wire [7:0] uio_oe,   // IOs: Bidirectional Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);


  //input wire clk,
  wire A8, A7, A6, A5, A4, A3, A2, A1;

assign uo_out[7:0] = {A8, A7, A6, A5, A4, A3, A2, A1};

assign uio_out = 8'b0;
reg clkA;

// use bidirectionals as outputs
    assign uio_oe = 8'b11111111;
    assign uio_out = 8'b0;
    
always @(posedge clk) begin
  if (!rst_n) begin
    clkA <= 0;
  end
  else begin
    clkA <= ~clkA;
  end
end

//Internal Wires
 wire [7:0] w_1;

//Instances os Modules
pulse_count_8_bits blk82_20 (
         .pulse (clkA),
         .counter (w_1)
     );

bus_to_wires blk28_22 (
         .out_2 (A3),
         .out_3 (A4),
         .out_1 (A2),
         .out_4 (A5),
         .out_0 (A1),
         .out_5 (A6),
         .out_7 (A8),
         .out_6 (A7),
         .in (w_1)
     );


endmodule
